netcdf columns_output_gfs_template {
dimensions:
        forecast_hour = unlimited ;
        sites = N_SITES ;
        height_bin = N_HEIGHT_BINS ;
        depth_bin = N_DEPTH_BINS ;
variables:
        float dlat(sites) ;
                dlat:long_name = "Desired site latitude" ;
                dlat:units = "degrees_north" ;
                dlat:_FillValue = 9.96921e+36f ;
        float dlon(sites) ;
                dlon:long_name = "Desired site longitude" ;
                dlon:units = "degrees_east" ;
                dlon:_FillValue = 9.96921e+36f ;
        string dsite(sites) ;
                dsite:long_name = "Desired site longname" ;
                dsite:units = "unitless" ;
        float mlat(sites) ;
                mlat:long_name = "Closest model grid point latitude" ;
                mlat:units = "degrees_north" ;
                mlat:_FillValue = 9.96921e+36f ;
        float mlon(sites) ;
                mlon:long_name = "Closest model grid point longitude" ;
                mlon:units = "degrees_east" ;
                mlon:_FillValue = 9.96921e+36f ;
        float distance(sites) ;
                distance:long_name = "Distance between desired and the model grid points" ;
                distance:units = "km" ;
                distance:_FillValue = 9.96921e+36f ;
        float height(height_bin) ;
                height:long_name = "Height" ;
                height:units = "m" ;
                height:positive = "up" ;
                height:description = "Heights are relative to ground level" ;
                height:_FillValue = 9.96921e+36f ;
        float depth(depth_bin) ;
                depth:long_name = "Depth" ;
                depth:units = "m" ;
                depth:positive = "down" ;
                depth:description = "Depths are relative to ground level" ;
                depth:_FillValue = 9.96921e+36f ;
        double model_initialization(forecast_hour) ;
                model_initialization:long_name = "Model initialization time" ;
                model_initialization:units = "seconds since 1970-01-01 00:00:00" ;
                model_initialization:_FillValue = 9.96921e+36 ;
        int forecast(forecast_hour) ;
                forecast:long_name = "Forecast hour" ;
                forecast:units = "hour" ;
                forecast:_FillValue = -9999 ;
        float p0(forecast_hour, sites, height_bin) ;
                p0:long_name = "Pressure at the closest model grid location" ;
                p0:units = "hPa" ;
                p0:_FillValue = 9.96921e+36f ;
        float p1(forecast_hour, sites, height_bin) ;
                p1:long_name = "Pressure calculated by bilinear interpolation via Scipy's griddata()" ;
                p1:units = "hPa" ;
                p1:_FillValue = 9.96921e+36f ;
        float t0(forecast_hour, sites, height_bin) ;
                t0:long_name = "Temperature at the closest model grid location" ;
                t0:units = "degC" ;
                t0:_FillValue = 9.96921e+36f ;
        float t1(forecast_hour, sites, height_bin) ;
                t1:long_name = "Temperature calculated by bilinear interpolation via Scipy's griddata()" ;
                t1:units = "degC" ;
                t1:_FillValue = 9.96921e+36f ;
        float qv0(forecast_hour, sites, height_bin) ;
                qv0:long_name = "Specific humidity at the closest model grid location" ;
                qv0:units = "g/kg" ;
                qv0:_FillValue = 9.96921e+36f ;
        float qv1(forecast_hour, sites, height_bin) ;
                qv1:long_name = "Specific humidity calculated by bilinear interpolation via Scipy's griddata()" ;
                qv1:units = "g/kg" ;
                qv1:_FillValue = 9.96921e+36f ;
        float r0(forecast_hour, sites, height_bin) ;
                r0:long_name = "Water vapor mixing ratio at the closest model grid location" ;
                r0:units = "g/kg" ;
                r0:_FillValue = 9.96921e+36f ;
        float r1(forecast_hour, sites, height_bin) ;
                r1:long_name = "Water vapor mixing ratio calculated by bilinear interpolation via Scipy's griddata()" ;
                r1:units = "g/kg" ;
                r1:_FillValue = 9.96921e+36f ;
        float tv0(forecast_hour, sites, height_bin) ;
                tv0:long_name = "Virtual temperature at the closest model grid location" ;
                tv0:units = "K" ;
                tv0:_FillValue = 9.96921e+36f ;
        float tv1(forecast_hour, sites, height_bin) ;
                tv1:long_name = "Virtual temperature calculated by bilinear interpolation via Scipy's griddata()" ;
                tv1:units = "K" ;
                tv1:_FillValue = 9.96921e+36f ;
        float lwc0(forecast_hour, sites, height_bin) ;
                lwc0:long_name = "Liquid water mixing ratio at the closest model grid location" ;
                lwc0:units = "kg/kg" ;
                lwc0:_FillValue = 9.96921e+36f ;
        float lwc1(forecast_hour, sites, height_bin) ;
                lwc1:long_name = "Liquid water mixing ratio calculated by bilinear interpolation via Scipy's griddata()" ;
                lwc1:units = "kg/kg" ;
                lwc1:_FillValue = 9.96921e+36f ;
        float totcc0(forecast_hour, sites, height_bin) ;
                totcc0:long_name = "Total cloud cover at the closest model grid location" ;
                totcc0:units = "%" ;
                totcc0:_FillValue = 9.96921e+36f ;
        float totcc1(forecast_hour, sites, height_bin) ;
                totcc1:long_name = "Total cloud cover calculated by bilinear interpolation via Scipy's griddata()" ;
                totcc1:units = "%" ;
                totcc1:_FillValue = 9.96921e+36f ;
        float wspd0(forecast_hour, sites, height_bin) ;
                wspd0:long_name = "Wind speed at the closest model grid location" ;
                wspd0:units = "m/s" ;
                wspd0:_FillValue = 9.96921e+36f ;
        float wspd1(forecast_hour, sites, height_bin) ;
                wspd1:long_name = "Wind speed calculated by bilinear interpolation via Scipy's griddata()" ;
                wspd1:units = "m/s" ;
                wspd1:_FillValue = 9.96921e+36f ;
        float u0(forecast_hour, sites, height_bin) ;
                u0:long_name = "u-component of wind at the closest model grid location" ;
                u0:units = "m/s" ;
                u0:_FillValue = 9.96921e+36f ;
        float u1(forecast_hour, sites, height_bin) ;
                u1:long_name = "u-component of wind calculated by bilinear interpolation via Scipy's griddata()" ;
                u1:units = "m/s" ;
                u1:_FillValue = 9.96921e+36f ;
        float v0(forecast_hour, sites, height_bin) ;
                v0:long_name = "v-component of wind at the closest model grid location" ;
                v0:units = "m/s" ;
                v0:_FillValue = 9.96921e+36f ;
        float v1(forecast_hour, sites, height_bin) ;
                v1:long_name = "v-component of wind calculated by bilinear interpolation via Scipy's griddata()" ;
                v1:units = "m/s" ;
                v1:_FillValue = 9.96921e+36f ;
        float w0(forecast_hour, sites, height_bin) ;
                w0:long_name = "w-component of wind at the closest model grid location" ;
                w0:units = "m/s" ;
                w0:_FillValue = 9.96921e+36f ;
        float w1(forecast_hour, sites, height_bin) ;
                w1:long_name = "w-component of wind calculated by bilinear interpolation via Scipy's griddata()" ;
                w1:units = "m/s" ;
                w1:_FillValue = 9.96921e+36f ;
        float soilt0(forecast_hour, sites, depth_bin) ;
                soilt0:long_name = "Soil temperature at the closest model grid location" ;
                soilt0:units = "K" ;
                soilt0:_FillValue = 9.96921e+36f ;
        float soilt1(forecast_hour, sites, depth_bin) ;
                soilt1:long_name = "Soil temperature calculated by bilinear interpolation via Scipy's griddata()" ;
                soilt1:units = "K" ;
                soilt1:_FillValue = 9.96921e+36f ;
        float soilm0(forecast_hour, sites, depth_bin) ;
                soilm0:long_name = "Volumetric soil moisture at the closest model grid location" ;
                soilm0:units = "Fraction" ;
                soilm0:_FillValue = 9.96921e+36f ;
        float soilm1(forecast_hour, sites, depth_bin) ;
                soilm1:long_name = "Volumetric soil moisture calculated by bilinear interpolation via Scipy's griddata()" ;
                soilm1:units = "Fraction" ;
                soilm1:_FillValue = 9.96921e+36f ;
        float pwv0(forecast_hour, sites) ;
                pwv0:long_name = "Precipitable water vapor at the closest model grid location" ;
                pwv0:units = "kg/m2" ;
                pwv0:_FillValue = 1.e+20f ;
        float pwv1(forecast_hour, sites) ;
                pwv1:long_name = "Precipitable water vapor calculated by bilinear interpolation via Scipy's griddata()" ;
                pwv1:units = "kg/m2" ;
                pwv1:_FillValue = 9.96921e+36f ;
        float pbl0(forecast_hour, sites) ;
                pbl0:long_name = "Planetary boundary layer height at the closest model grid location" ;
                pbl0:units = "m" ;
                pbl0:_FillValue = 1.e+20f ;
        float pbl1(forecast_hour, sites) ;
                pbl1:long_name = "Planetary boundary layer height calculated by bilinear interpolation via Scipy's griddata()" ;
                pbl1:units = "m" ;
                pbl1:_FillValue = 9.96921e+36f ;
        float stemp0(forecast_hour, sites) ;
                stemp0:long_name = "Surface skin temperature at the closest model grid location" ;
                stemp0:units = "degC" ;
                stemp0:_FillValue = 1.e+20f ;
        float stemp1(forecast_hour, sites) ;
                stemp1:long_name = "Surface skin temperature calculated by bilinear interpolation via Scipy's griddata()" ;
                stemp1:units = "degC" ;
                stemp1:_FillValue = 9.96921e+36f ;
        float lflux0(forecast_hour, sites) ;
                lflux0:long_name = "Latent heat flux at the closest model grid location" ;
                lflux0:description = "Averaged over previous N forecast hours" ;
                lflux0:units = "W/m2" ;
                lflux0:_FillValue = 1.e+20f ;
        float lflux1(forecast_hour, sites) ;
                lflux1:long_name = "Latent heat flux calculated by bilinear interpolation via Scipy's griddata()" ;
                lflux1:description = "Averaged over previous N forecast hours" ;
                lflux1:units = "W/m2" ;
                lflux1:_FillValue = 9.96921e+36f ;
        float sflux0(forecast_hour, sites) ;
                sflux0:long_name = "Sensible heat flux at the closest model grid location" ;
                sflux0:description = "Averaged over previous N forecast hours" ;
                sflux0:units = "W/m2" ;
                sflux0:_FillValue = 1.e+20f ;
        float sflux1(forecast_hour, sites) ;
                sflux1:long_name = "Sensible heat flux calculated by bilinear interpolation via Scipy's griddata()" ;
                sflux1:description = "Averaged over previous N forecast hours" ;
                sflux1:units = "W/m2" ;
                sflux1:_FillValue = 9.96921e+36f ;
        float gflux0(forecast_hour, sites) ;
                gflux0:long_name = "Ground heat flux at the closest model grid location" ;
                gflux0:description = "Averaged over previous N forecast hours" ;
                gflux0:units = "W/m2" ;
                gflux0:_FillValue = 1.e+20f ;
        float gflux1(forecast_hour, sites) ;
                gflux1:long_name = "Ground heat flux calculated by bilinear interpolation via Scipy's griddata()" ;
                gflux1:description = "Averaged over previous N forecast hours" ;
                gflux1:units = "W/m2" ;
                gflux1:_FillValue = 9.96921e+36f ;
        float dswsfc0(forecast_hour, sites) ;
                dswsfc0:long_name = "Downwelling SW flux at the surface at the closest model grid location" ;
                dswsfc0:description = "Averaged over previous N forecast hours" ;
                dswsfc0:units = "W/m2" ;
                dswsfc0:_FillValue = 1.e+20f ;
        float dswsfc1(forecast_hour, sites) ;
                dswsfc1:long_name = "Downwelling SW flux at the surface calculated by bilinear interpolation via Scipy's griddata()" ;
                dswsfc1:description = "Averaged over previous N forecast hours" ;
                dswsfc1:units = "W/m2" ;
                dswsfc1:_FillValue = 9.96921e+36f ;
        float uswsfc0(forecast_hour, sites) ;
                uswsfc0:long_name = "Upwelling SW flux at the surface at the closest model grid location" ;
                uswsfc0:description = "Averaged over previous N forecast hours" ;
                uswsfc0:units = "W/m2" ;
                uswsfc0:_FillValue = 1.e+20f ;
        float uswsfc1(forecast_hour, sites) ;
                uswsfc1:long_name = "Upwelling SW flux at the surface calculated by bilinear interpolation via Scipy's griddata()" ;
                uswsfc1:description = "Averaged over previous N forecast hours" ;
                uswsfc1:units = "W/m2" ;
                uswsfc1:_FillValue = 9.96921e+36f ;
        float uswtoa0(forecast_hour, sites) ;
                uswtoa0:long_name = "Upwelling shortwave flux at the top of atmosphere at the closest model grid location" ;
                uswtoa0:description = "Averaged over previous N forecast hours" ;
                uswtoa0:units = "W/m2" ;
                uswtoa0:_FillValue = 9.96921e+36f ;
        float uswtoa1(forecast_hour, sites) ;
                uswtoa1:long_name = "Upwelling shortwave flux at the top of atmosphere calculated by bilinear interpolation via Scipy's griddata()" ;
                uswtoa1:description = "Averaged over previous N forecast hours" ;
                uswtoa1:units = "W/m2" ;
                uswtoa1:_FillValue = 9.96921e+36f ;
        float ulwtoa0(forecast_hour, sites) ;
                ulwtoa0:long_name = "Upwelling LW flux at the TOA at the closest model grid location" ;
                ulwtoa0:description = "Averaged over previous N forecast hours" ;
                ulwtoa0:units = "W/m2" ;
                ulwtoa0:_FillValue = 1.e+20f ;
        float ulwtoa1(forecast_hour, sites) ;
                ulwtoa1:long_name = "Upwelling LW flux at the TOA calculated by bilinear interpolation via Scipy's griddata()" ;
                ulwtoa1:description = "Averaged over previous N forecast hours" ;
                ulwtoa1:units = "W/m2" ;
                ulwtoa1:_FillValue = 9.96921e+36f ;
        float dlwsfc0(forecast_hour, sites) ;
                dlwsfc0:long_name = "Downwelling LW flux at the surface at the closest model grid location" ;
                dlwsfc0:description = "Averaged over previous N forecast hours" ;
                dlwsfc0:units = "W/m2" ;
                dlwsfc0:_FillValue = 1.e+20f ;
        float dlwsfc1(forecast_hour, sites) ;
                dlwsfc1:long_name = "Downwelling LW flux at the surface calculated by bilinear interpolation via Scipy's griddata()" ;
                dlwsfc1:description = "Averaged over previous N forecast hours" ;
                dlwsfc1:units = "W/m2" ;
                dlwsfc1:_FillValue = 9.96921e+36f ;
        float ulwsfc0(forecast_hour, sites) ;
                ulwsfc0:long_name = "Upwelling LW flux at the surface at the closest model grid location" ;
                ulwsfc0:description = "Averaged over previous N forecast hours" ;
                ulwsfc0:units = "W/m2" ;
                ulwsfc0:_FillValue = 1.e+20f ;
        float ulwsfc1(forecast_hour, sites) ;
                ulwsfc1:long_name = "Upwelling LW flux at the surface calculated by bilinear interpolation via Scipy's griddata()" ;
                ulwsfc1:description = "Averaged over previous N forecast hours" ;
                ulwsfc1:units = "W/m2" ;
                ulwsfc1:_FillValue = 9.96921e+36f ;
        float tcc0(forecast_hour, sites) ;
                tcc0:long_name = "Total cloud cover fraction at the closest model grid location" ;
                tcc0:units = "%" ;
                tcc0:_FillValue = 1.e+20f ;
        float tcc1(forecast_hour, sites) ;
                tcc1:long_name = "Total cloud cover fraction calculated by bilinear interpolation via Scipy's griddata()" ;
                tcc1:units = "%" ;
                tcc1:_FillValue = 9.96921e+36f ;
        float lcc0(forecast_hour, sites) ;
                lcc0:long_name = "Low cloud cover fraction at the closest model grid location" ;
                lcc0:units = "%" ;
                lcc0:_FillValue = 1.e+20f ;
        float lcc1(forecast_hour, sites) ;
                lcc1:long_name = "Low cloud cover fraction calculated by bilinear interpolation via Scipy's griddata()" ;
                lcc1:units = "%" ;
                lcc1:_FillValue = 9.96921e+36f ;
        float mcc0(forecast_hour, sites) ;
                mcc0:long_name = "Medium cloud cover fraction at the closest model grid location" ;
                mcc0:units = "%" ;
                mcc0:_FillValue = 1.e+20f ;
        float mcc1(forecast_hour, sites) ;
                mcc1:long_name = "Medium cloud cover fraction calculated by bilinear interpolation via Scipy's griddata()" ;
                mcc1:units = "%" ;
                mcc1:_FillValue = 9.96921e+36f ;
        float hcc0(forecast_hour, sites) ;
                hcc0:long_name = "High cloud cover fraction at the closest model grid location" ;
                hcc0:units = "%" ;
                hcc0:_FillValue = 1.e+20f ;
        float hcc1(forecast_hour, sites) ;
                hcc1:long_name = "High cloud cover fraction calculated by bilinear interpolation via Scipy's griddata()" ;
                hcc1:units = "%" ;
                hcc1:_FillValue = 9.96921e+36f ;
        float vis0(forecast_hour, sites) ;
                vis0:long_name = "Visibility at the closest model grid location" ;
                vis0:units = "m" ;
                vis0:_FillValue = 1.e+20f ;
        float vis1(forecast_hour, sites) ;
                vis1:long_name = "Visibility calculated by bilinear interpolation via Scipy's griddata()" ;
                vis1:units = "m" ;
                vis1:_FillValue = 9.96921e+36f ;
        float crefl0(forecast_hour, sites) ;
                crefl0:long_name = "Composite reflectivity at the closest model grid location" ;
                crefl0:units = "dBZ" ;
                crefl0:_FillValue = 1.e+20f ;
        float crefl1(forecast_hour, sites) ;
                crefl1:long_name = "Composite reflectivity calculated by bilinear interpolation via Scipy's griddata()" ;
                crefl1:units = "dBZ" ;
                crefl1:_FillValue = 9.96921e+36f ;
        float terr0(forecast_hour, sites) ;
                terr0:long_name = "Terrain height at the closest model grid location" ;
                terr0:units = "m" ;
                terr0:_FillValue = 1.e+20f ;
        float terr1(forecast_hour, sites) ;
                terr1:long_name = "Terrain height calculated by bilinear interpolation via Scipy's griddata()" ;
                terr1:units = "m" ;
                terr1:_FillValue = 9.96921e+36f ;
        float ustar0(forecast_hour, sites) ;
                ustar0:long_name = "Friction velocity at the closest model grid location" ;
                ustar0:units = "m/s" ;
                ustar0:_FillValue = 9.96921e+36f ;
        float ustar1(forecast_hour, sites) ;
                ustar1:long_name = "Friction velocity calculated by bilinear interpolation via Scipy's griddata()" ;
                ustar1:units = "m/s" ;
                ustar1:_FillValue = 9.96921e+36f ;
        float prate0(forecast_hour, sites) ;
                prate0:long_name = "Precipitation rate at the closest model grid location" ;
                prate0:units = "kg/m2s" ;
                prate0:_FillValue = 9.96921e+36f ;
        float prate1(forecast_hour, sites) ;
                prate1:long_name = "Precipitation rate calculated by bilinear interpolation via Scipy's griddata()" ;
                prate1:units = "kg/m2s" ;
                prate1:_FillValue = 9.96921e+36f ;
        float csnow0(forecast_hour, sites) ;
                csnow0:long_name = "Categorical snow at the closest model grid location (1-yes, 0-no)" ;
                csnow0:units = "unitless" ;
                csnow0:_FillValue = 9.96921e+36f ;
        float csnow1(forecast_hour, sites) ;
                csnow1:long_name = "Categorical snow at the closest model grid location (1-yes, 0-no)" ;
                csnow1:units = "unitless" ;
                csnow1:_FillValue = 9.96921e+36f ;
        float psfc0(forecast_hour, sites) ;
                psfc0:long_name = "Pressure at the surface at the closest model grid location" ;
                psfc0:units = "hPa" ;
                psfc0:_FillValue = 1.e+20f ;
        float psfc1(forecast_hour, sites) ;
                psfc1:long_name = "Pressure at the surface calculated by bilinear interpolation via Scipy's griddata()" ;
                psfc1:units = "hPa" ;
                psfc1:_FillValue = 9.96921e+36f ;
        float tsfc0(forecast_hour, sites) ;
                tsfc0:long_name = "Temperature at 2-m at the closest model grid location" ;
                tsfc0:units = "degC" ;
                tsfc0:_FillValue = 1.e+20f ;
        float tsfc1(forecast_hour, sites) ;
                tsfc1:long_name = "Temperature at 2-m calculated by bilinear interpolation via Scipy's griddata()" ;
                tsfc1:units = "degC" ;
                tsfc1:_FillValue = 9.96921e+36f ;
        float dpsfc0(forecast_hour, sites) ;
                dpsfc0:long_name = "Dew point temperature at 2-m at the closest model grid location" ;
                dpsfc0:units = "degC" ;
                dpsfc0:_FillValue = 1.e+20f ;
        float dpsfc1(forecast_hour, sites) ;
                dpsfc1:long_name = "Dew point temperature at 2-m calculated by bilinear interpolation via Scipy's griddata()" ;
                dpsfc1:units = "degC" ;
                dpsfc1:_FillValue = 9.96921e+36f ;
        float rhsfc0(forecast_hour, sites) ;
                rhsfc0:long_name = "Relative humidity at 2-m at the closest model grid location" ;
                rhsfc0:units = "%" ;
                rhsfc0:_FillValue = 9.96921e+36f ;
        float rhsfc1(forecast_hour, sites) ;
                rhsfc1:long_name = "Relative humidity at 2-m calculated by bilinear interpolation via Scipy's griddata()" ;
                rhsfc1:units = "%" ;
                rhsfc1:_FillValue = 9.96921e+36f ;
        float qvsfc0(forecast_hour, sites) ;
                qvsfc0:long_name = "Specific humidity at 2-m at the closest model grid location" ;
                qvsfc0:units = "g/kg" ;
                qvsfc0:_FillValue = 1.e+20f ;
        float qvsfc1(forecast_hour, sites) ;
                qvsfc1:long_name = "Specific humidity at 2-m calculated by bilinear interpolation via Scipy's griddata()" ;
                qvsfc1:units = "g/kg" ;
                qvsfc1:_FillValue = 9.96921e+36f ;
        float rsfc0(forecast_hour, sites) ;
                rsfc0:long_name = "Water vapor mixing ratio at 2-m at the closest model grid location" ;
                rsfc0:units = "g/kg" ;
                rsfc0:_FillValue = 9.96921e+36f ;
        float rsfc1(forecast_hour, sites) ;
                rsfc1:long_name = "Water vapor mixing ratio at 2-m calculated by bilinear interpolation via Scipy's griddata()" ;
                rsfc1:units = "g/kg" ;
                rsfc1:_FillValue = 9.96921e+36f ;
        float usfc0(forecast_hour, sites) ;
                usfc0:long_name = "U-component of wind at 10-m at the closest model grid location" ;
                usfc0:units = "m/s" ;
                usfc0:_FillValue = 1.e+20f ;
        float usfc1(forecast_hour, sites) ;
                usfc1:long_name = "U-component of wind at 10-m calculated by bilinear interpolation via Scipy's griddata()" ;
                usfc1:units = "m/s" ;
                usfc1:_FillValue = 9.96921e+36f ;
        float vsfc0(forecast_hour, sites) ;
                vsfc0:long_name = "V-component of wind at 10-m at the closest model grid location" ;
                vsfc0:units = "m/s" ;
                vsfc0:_FillValue = 1.e+20f ;
        float vsfc1(forecast_hour, sites) ;
                vsfc1:long_name = "V-component of wind at 10-m calculated by bilinear interpolation via Scipy's griddata()" ;
                vsfc1:units = "m/s" ;
                vsfc1:_FillValue = 9.96921e+36f ;
        float u80m0(forecast_hour, sites) ;
                u80m0:long_name = "U-component of wind at 80-m at the closest model grid location" ;
                u80m0:units = "m/s" ;
                u80m0:_FillValue = 9.96921e+36f ;
        float u80m1(forecast_hour, sites) ;
                u80m1:long_name = "U-component of wind at 80-m calculated by bilinear interpolation via Scipy's griddata()" ;
                u80m1:units = "m/s" ;
                u80m1:_FillValue = 9.96921e+36f ;
        float v80m0(forecast_hour, sites) ;
                v80m0:long_name = "V-component of wind at 80-m at the closest model grid location" ;
                v80m0:units = "m/s" ;
                v80m0:_FillValue = 9.96921e+36f ;
        float v80m1(forecast_hour, sites) ;
                v80m1:long_name = "V-component of wind at 80-m calculated by bilinear interpolation via Scipy's griddata()" ;
                v80m1:units = "m/s" ;
                v80m1:_FillValue = 9.96921e+36f ;

// global attributes:
                :title = "Vertical profiles / point values at profiling sites of interest" ;
                :institution = "NOAA Global Systems Laboratory (GSL)" ;
                :contact = "dsg.its.gsl@noaa.gov, dave.turner@noaa.gov" ;
                :source = SOURCE_FILE ;
                :model = "GFS V16 (0.25deg)" ;
	        :model_initialization = MODEL_INIT ;
                :version = CODE_VERSION ;
                :references = "https://github.com/NOAA-GSL/column-extractor" ;
                :Conventions = "CF-1.10" ;
                :date_file_created = FILE_CREATION_TIME ;
}
